library verilog;
use verilog.vl_types.all;
entity contador_assincrono_ffjk_vlg_vec_tst is
end contador_assincrono_ffjk_vlg_vec_tst;
